library ieee;
use ieee.std_logic_1164.all;
use work.float_pkg.all;
--use work.myTypes.all;
use work.fixed_pkg.all;
use work.float_pkg.all;

package LUT is
  	constant LIMIT_1 : float16 := to_float(0.5, 5, 10);
  	constant LIMIT_2 : float16 := to_float(1.0, 5, 10);
  	constant LIMIT_3 : float16 := to_float(1.5, 5, 10);
  	constant LIMIT_4 : float16 := to_float(2.0, 5, 10);
  	constant N_1: integer := 128;
  	constant N_2: integer := 64;
  	constant N_3: integer := 32;
	constant N_4: integer := 32;
    	constant LUT_SIZE : integer := N_1 + N_2 +N_3 + N_4;

    	type lut_array is array (0 to LUT_SIZE-1) of float16;

    constant lut_values : lut_array := (


x"3800", --   0  (x=0.0000, sig=0.500000)
x"3808", --   1  (x=0.0039, sig=0.503906)
x"3810", --   2  (x=0.0078, sig=0.507812)
x"3818", --   3  (x=0.0117, sig=0.511719)
x"3820", --   4  (x=0.0156, sig=0.515625)
x"3828", --   5  (x=0.0195, sig=0.519531)
x"3830", --   6  (x=0.0234, sig=0.523438)
x"3838", --   7  (x=0.0273, sig=0.527344)
x"3840", --   8  (x=0.0312, sig=0.531250)
x"3848", --   9  (x=0.0352, sig=0.535156)
x"3850", --  10  (x=0.0391, sig=0.539062)
x"3858", --  11  (x=0.0430, sig=0.542969)
x"3860", --  12  (x=0.0469, sig=0.546875)
x"3868", --  13  (x=0.0508, sig=0.550781)
x"386f", --  14  (x=0.0547, sig=0.554199)
x"3877", --  15  (x=0.0586, sig=0.558105)
x"387f", --  16  (x=0.0625, sig=0.562012)
x"3887", --  17  (x=0.0664, sig=0.565918)
x"388f", --  18  (x=0.0703, sig=0.569824)
x"3897", --  19  (x=0.0742, sig=0.573730)
x"389f", --  20  (x=0.0781, sig=0.577637)
x"38a6", --  21  (x=0.0820, sig=0.581055)
x"38ae", --  22  (x=0.0859, sig=0.584961)
x"38b6", --  23  (x=0.0898, sig=0.588867)
x"38be", --  24  (x=0.0938, sig=0.592773)
x"38c5", --  25  (x=0.0977, sig=0.596191)
x"38cd", --  26  (x=0.1016, sig=0.600098)
x"38d5", --  27  (x=0.1055, sig=0.604004)
x"38dd", --  28  (x=0.1094, sig=0.607910)
x"38e4", --  29  (x=0.1133, sig=0.611328)
x"38ec", --  30  (x=0.1172, sig=0.615234)
x"38f3", --  31  (x=0.1211, sig=0.618652)
x"38fb", --  32  (x=0.1250, sig=0.622559)
x"3902", --  33  (x=0.1289, sig=0.625977)
x"390a", --  34  (x=0.1328, sig=0.629883)
x"3912", --  35  (x=0.1367, sig=0.633789)
x"3918", --  36  (x=0.1406, sig=0.636719)
x"3920", --  37  (x=0.1445, sig=0.640625)
x"3927", --  38  (x=0.1484, sig=0.644043)
x"392f", --  39  (x=0.1523, sig=0.647949)
x"3936", --  40  (x=0.1562, sig=0.651367)
x"393d", --  41  (x=0.1602, sig=0.654785)
x"3945", --  42  (x=0.1641, sig=0.658691)
x"394c", --  43  (x=0.1680, sig=0.662109)
x"3953", --  44  (x=0.1719, sig=0.665527)
x"395a", --  45  (x=0.1758, sig=0.668945)
x"3961", --  46  (x=0.1797, sig=0.672363)
x"3968", --  47  (x=0.1836, sig=0.675781)
x"396f", --  48  (x=0.1875, sig=0.679199)
x"3976", --  49  (x=0.1914, sig=0.682617)
x"397d", --  50  (x=0.1953, sig=0.686035)
x"3983", --  51  (x=0.1992, sig=0.688965)
x"398b", --  52  (x=0.2031, sig=0.692871)
x"3992", --  53  (x=0.2070, sig=0.696289)
x"3998", --  54  (x=0.2109, sig=0.699219)
x"399e", --  55  (x=0.2148, sig=0.702148)
x"39a5", --  56  (x=0.2188, sig=0.705566)
x"39ac", --  57  (x=0.2227, sig=0.708984)
x"39b2", --  58  (x=0.2266, sig=0.711914)
x"39ba", --  59  (x=0.2305, sig=0.715820)
x"39c0", --  60  (x=0.2344, sig=0.718750)
x"39c6", --  61  (x=0.2383, sig=0.721680)
x"39cc", --  62  (x=0.2422, sig=0.724609)
x"39d3", --  63  (x=0.2461, sig=0.728027)
x"39d9", --  64  (x=0.2500, sig=0.730957)
x"39df", --  65  (x=0.2539, sig=0.733887)
x"39e6", --  66  (x=0.2578, sig=0.737305)
x"39eb", --  67  (x=0.2617, sig=0.739746)
x"39f2", --  68  (x=0.2656, sig=0.743164)
x"39f9", --  69  (x=0.2695, sig=0.746582)
x"39fe", --  70  (x=0.2734, sig=0.749023)
x"3a04", --  71  (x=0.2773, sig=0.751953)
x"3a0b", --  72  (x=0.2812, sig=0.755371)
x"3a10", --  73  (x=0.2852, sig=0.757812)
x"3a16", --  74  (x=0.2891, sig=0.760742)
x"3a1c", --  75  (x=0.2930, sig=0.763672)
x"3a22", --  76  (x=0.2969, sig=0.766602)
x"3a26", --  77  (x=0.3008, sig=0.768555)
x"3a2c", --  78  (x=0.3047, sig=0.771484)
x"3a32", --  79  (x=0.3086, sig=0.774414)
x"3a37", --  80  (x=0.3125, sig=0.776855)
x"3a3d", --  81  (x=0.3164, sig=0.779785)
x"3a43", --  82  (x=0.3203, sig=0.782715)
x"3a48", --  83  (x=0.3242, sig=0.785156)
x"3a4d", --  84  (x=0.3281, sig=0.787598)
x"3a53", --  85  (x=0.3320, sig=0.790527)
x"3a58", --  86  (x=0.3359, sig=0.792969)
x"3a5d", --  87  (x=0.3398, sig=0.795410)
x"3a63", --  88  (x=0.3438, sig=0.798340)
x"3a68", --  89  (x=0.3477, sig=0.800781)
x"3a6d", --  90  (x=0.3516, sig=0.803223)
x"3a72", --  91  (x=0.3555, sig=0.805664)
x"3a77", --  92  (x=0.3594, sig=0.808105)
x"3a7b", --  93  (x=0.3633, sig=0.810059)
x"3a80", --  94  (x=0.3672, sig=0.812500)
x"3a86", --  95  (x=0.3711, sig=0.815430)
x"3a8b", --  96  (x=0.3750, sig=0.817871)
x"3a8f", --  97  (x=0.3789, sig=0.819824)
x"3a93", --  98  (x=0.3828, sig=0.821777)
x"3a99", --  99  (x=0.3867, sig=0.824707)
x"3a9d", -- 100  (x=0.3906, sig=0.826660)
x"3aa2", -- 101  (x=0.3945, sig=0.829102)
x"3aa6", -- 102  (x=0.3984, sig=0.831055)
x"3aaa", -- 103  (x=0.4023, sig=0.833008)
x"3aaf", -- 104  (x=0.4062, sig=0.835449)
x"3ab4", -- 105  (x=0.4102, sig=0.837891)
x"3ab8", -- 106  (x=0.4141, sig=0.839844)
x"3abd", -- 107  (x=0.4180, sig=0.842285)
x"3ac1", -- 108  (x=0.4219, sig=0.844238)
x"3ac5", -- 109  (x=0.4258, sig=0.846191)
x"3ac8", -- 110  (x=0.4297, sig=0.847656)
x"3acc", -- 111  (x=0.4336, sig=0.849609)
x"3ad1", -- 112  (x=0.4375, sig=0.852051)
x"3ad5", -- 113  (x=0.4414, sig=0.854004)
x"3ad9", -- 114  (x=0.4453, sig=0.855957)
x"3adc", -- 115  (x=0.4492, sig=0.857422)
x"3ae1", -- 116  (x=0.4531, sig=0.859863)
x"3ae4", -- 117  (x=0.4570, sig=0.861328)
x"3ae8", -- 118  (x=0.4609, sig=0.863281)
x"3aeb", -- 119  (x=0.4648, sig=0.864746)
x"3af0", -- 120  (x=0.4688, sig=0.867188)
x"3af3", -- 121  (x=0.4727, sig=0.868652)
x"3af7", -- 122  (x=0.4766, sig=0.870605)
x"3afa", -- 123  (x=0.4805, sig=0.872070)
x"3afd", -- 124  (x=0.4844, sig=0.873535)
x"3b02", -- 125  (x=0.4883, sig=0.875977)
x"3b05", -- 126  (x=0.4922, sig=0.877441)
x"3b08", -- 127  (x=0.4961, sig=0.878906)
x"3b0b", -- 128  (x=0.5000, sig=0.880371)
x"3b13", -- 129  (x=0.5078, sig=0.884277)
x"3b19", -- 130  (x=0.5156, sig=0.887207)
x"3b20", -- 131  (x=0.5234, sig=0.890625)
x"3b26", -- 132  (x=0.5312, sig=0.893555)
x"3b2b", -- 133  (x=0.5391, sig=0.895996)
x"3b31", -- 134  (x=0.5469, sig=0.898926)
x"3b38", -- 135  (x=0.5547, sig=0.902344)
x"3b3d", -- 136  (x=0.5625, sig=0.904785)
x"3b42", -- 137  (x=0.5703, sig=0.907227)
x"3b48", -- 138  (x=0.5781, sig=0.910156)
x"3b4d", -- 139  (x=0.5859, sig=0.912598)
x"3b52", -- 140  (x=0.5938, sig=0.915039)
x"3b57", -- 141  (x=0.6016, sig=0.917480)
x"3b5b", -- 142  (x=0.6094, sig=0.919434)
x"3b60", -- 143  (x=0.6172, sig=0.921875)
x"3b65", -- 144  (x=0.6250, sig=0.924316)
x"3b68", -- 145  (x=0.6328, sig=0.925781)
x"3b6d", -- 146  (x=0.6406, sig=0.928223)
x"3b71", -- 147  (x=0.6484, sig=0.930176)
x"3b76", -- 148  (x=0.6562, sig=0.932617)
x"3b79", -- 149  (x=0.6641, sig=0.934082)
x"3b7d", -- 150  (x=0.6719, sig=0.936035)
x"3b80", -- 151  (x=0.6797, sig=0.937500)
x"3b86", -- 152  (x=0.6875, sig=0.940430)
x"3b89", -- 153  (x=0.6953, sig=0.941895)
x"3b8b", -- 154  (x=0.7031, sig=0.942871)
x"3b8f", -- 155  (x=0.7109, sig=0.944824)
x"3b92", -- 156  (x=0.7188, sig=0.946289)
x"3b96", -- 157  (x=0.7266, sig=0.948242)
x"3b99", -- 158  (x=0.7344, sig=0.949707)
x"3b9b", -- 159  (x=0.7422, sig=0.950684)
x"3b9f", -- 160  (x=0.7500, sig=0.952637)
x"3ba2", -- 161  (x=0.7578, sig=0.954102)
x"3ba4", -- 162  (x=0.7656, sig=0.955078)
x"3ba8", -- 163  (x=0.7734, sig=0.957031)
x"3baa", -- 164  (x=0.7812, sig=0.958008)
x"3bac", -- 165  (x=0.7891, sig=0.958984)
x"3baf", -- 166  (x=0.7969, sig=0.960449)
x"3bb1", -- 167  (x=0.8047, sig=0.961426)
x"3bb3", -- 168  (x=0.8125, sig=0.962402)
x"3bb7", -- 169  (x=0.8203, sig=0.964355)
x"3bb9", -- 170  (x=0.8281, sig=0.965332)
x"3bba", -- 171  (x=0.8359, sig=0.965820)
x"3bbc", -- 172  (x=0.8438, sig=0.966797)
x"3bbe", -- 173  (x=0.8516, sig=0.967773)
x"3bc0", -- 174  (x=0.8594, sig=0.968750)
x"3bc2", -- 175  (x=0.8672, sig=0.969727)
x"3bc4", -- 176  (x=0.8750, sig=0.970703)
x"3bc6", -- 177  (x=0.8828, sig=0.971680)
x"3bc8", -- 178  (x=0.8906, sig=0.972656)
x"3bc9", -- 179  (x=0.8984, sig=0.973145)
x"3bcb", -- 180  (x=0.9062, sig=0.974121)
x"3bcd", -- 181  (x=0.9141, sig=0.975098)
x"3bcd", -- 182  (x=0.9219, sig=0.975098)
x"3bcf", -- 183  (x=0.9297, sig=0.976074)
x"3bd1", -- 184  (x=0.9375, sig=0.977051)
x"3bd3", -- 185  (x=0.9453, sig=0.978027)
x"3bd3", -- 186  (x=0.9531, sig=0.978027)
x"3bd5", -- 187  (x=0.9609, sig=0.979004)
x"3bd7", -- 188  (x=0.9688, sig=0.979980)
x"3bd7", -- 189  (x=0.9766, sig=0.979980)
x"3bd9", -- 190  (x=0.9844, sig=0.980957)
x"3bdb", -- 191  (x=0.9922, sig=0.981934)
x"3bdb", -- 192  (x=1.0000, sig=0.981934)
x"3bdd", -- 193  (x=1.0156, sig=0.982910)
x"3bdf", -- 194  (x=1.0312, sig=0.983887)
x"3be0", -- 195  (x=1.0469, sig=0.984375)
x"3be2", -- 196  (x=1.0625, sig=0.985352)
x"3be4", -- 197  (x=1.0781, sig=0.986328)
x"3be6", -- 198  (x=1.0938, sig=0.987305)
x"3be8", -- 199  (x=1.1094, sig=0.988281)
x"3bea", -- 200  (x=1.1250, sig=0.989258)
x"3bea", -- 201  (x=1.1406, sig=0.989258)
x"3bec", -- 202  (x=1.1562, sig=0.990234)
x"3bee", -- 203  (x=1.1719, sig=0.991211)
x"3bee", -- 204  (x=1.1875, sig=0.991211)
x"3bf0", -- 205  (x=1.2031, sig=0.992188)
x"3bf0", -- 206  (x=1.2188, sig=0.992188)
x"3bf2", -- 207  (x=1.2344, sig=0.993164)
x"3bf2", -- 208  (x=1.2500, sig=0.993164)
x"3bf4", -- 209  (x=1.2656, sig=0.994141)
x"3bf4", -- 210  (x=1.2812, sig=0.994141)
x"3bf4", -- 211  (x=1.2969, sig=0.994141)
x"3bf6", -- 212  (x=1.3125, sig=0.995117)
x"3bf6", -- 213  (x=1.3281, sig=0.995117)
x"3bf6", -- 214  (x=1.3438, sig=0.995117)
x"3bf8", -- 215  (x=1.3594, sig=0.996094)
x"3bf8", -- 216  (x=1.3750, sig=0.996094)
x"3bf8", -- 217  (x=1.3906, sig=0.996094)
x"3bf8", -- 218  (x=1.4062, sig=0.996094)
x"3bfa", -- 219  (x=1.4219, sig=0.997070)
x"3bfa", -- 220  (x=1.4375, sig=0.997070)
x"3bfa", -- 221  (x=1.4531, sig=0.997070)
x"3bfa", -- 222  (x=1.4688, sig=0.997070)
x"3bfa", -- 223  (x=1.4844, sig=0.997070)
x"3bfa", -- 224  (x=1.5000, sig=0.997070)
x"3bfc", -- 225  (x=1.5166, sig=0.998047)
x"3bfc", -- 226  (x=1.5322, sig=0.998047)
x"3bfc", -- 227  (x=1.5488, sig=0.998047)
x"3bfc", -- 228  (x=1.5645, sig=0.998047)
x"3bfc", -- 229  (x=1.5811, sig=0.998047)
x"3bfc", -- 230  (x=1.5967, sig=0.998047)
x"3bfc", -- 231  (x=1.6133, sig=0.998047)
x"3bfc", -- 232  (x=1.6289, sig=0.998047)
x"3bfe", -- 233  (x=1.6455, sig=0.999023)
x"3bfe", -- 234  (x=1.6611, sig=0.999023)
x"3bfe", -- 235  (x=1.6777, sig=0.999023)
x"3bfe", -- 236  (x=1.6934, sig=0.999023)
x"3bfe", -- 237  (x=1.7100, sig=0.999023)
x"3bfe", -- 238  (x=1.7256, sig=0.999023)
x"3bfe", -- 239  (x=1.7422, sig=0.999023)
x"3bfe", -- 240  (x=1.7578, sig=0.999023)
x"3bfe", -- 241  (x=1.7744, sig=0.999023)
x"3bfe", -- 242  (x=1.7900, sig=0.999023)
x"3bfe", -- 243  (x=1.8066, sig=0.999023)
x"3bfe", -- 244  (x=1.8223, sig=0.999023)
x"3bfe", -- 245  (x=1.8389, sig=0.999023)
x"3bfe", -- 246  (x=1.8545, sig=0.999023)
x"3bfe", -- 247  (x=1.8711, sig=0.999023)
x"3bfe", -- 248  (x=1.8867, sig=0.999023)
x"3bfe", -- 249  (x=1.9033, sig=0.999023)
x"3c00", -- 250  (x=1.9199, sig=1.000000)
x"3c00", -- 251  (x=1.9355, sig=1.000000)
x"3c00", -- 252  (x=1.9512, sig=1.000000)
x"3c00", -- 253  (x=1.9678, sig=1.000000)
x"3c00", -- 254  (x=1.9844, sig=1.000000)
x"3c00" -- 255  (x=2.0000, sig=1.000000)




    );
end package LUT;

