library ieee;
use ieee.std_logic_1164.all;
use work.float_pkg.all;
--use work.myTypes.all;
use work.fixed_pkg.all;
use work.float_pkg.all;

package LUT is
  	constant LIMIT_1 : float16 := to_float(0.5, 5, 10);
  	constant LIMIT_2 : float16 := to_float(1.0, 5, 10);
  	constant LIMIT_3 : float16 := to_float(1.5, 5, 10);
  	constant LIMIT_4 : float16 := to_float(2.0, 5, 10);
  	constant N_1: integer := 256;
  	constant N_2: integer := 128;
  	constant N_3: integer := 64;
	constant N_4: integer := 64;
    	constant LUT_SIZE : integer := N_1 + N_2 +N_3 + N_4;

    	type lut_array is array (0 to LUT_SIZE-1) of float16;

    constant lut_values : lut_array := (
x"3800", --   0  (x=0.0000, sig=0.500000)
x"3804", --   1  (x=0.0020, sig=0.501953)
x"3808", --   2  (x=0.0039, sig=0.503906)
x"380c", --   3  (x=0.0059, sig=0.505859)
x"3810", --   4  (x=0.0078, sig=0.507812)
x"3814", --   5  (x=0.0098, sig=0.509766)
x"3818", --   6  (x=0.0117, sig=0.511719)
x"381c", --   7  (x=0.0137, sig=0.513672)
x"3820", --   8  (x=0.0156, sig=0.515625)
x"3824", --   9  (x=0.0176, sig=0.517578)
x"3828", --  10  (x=0.0195, sig=0.519531)
x"382c", --  11  (x=0.0215, sig=0.521484)
x"3830", --  12  (x=0.0234, sig=0.523438)
x"3834", --  13  (x=0.0254, sig=0.525391)
x"3838", --  14  (x=0.0273, sig=0.527344)
x"383c", --  15  (x=0.0293, sig=0.529297)
x"3840", --  16  (x=0.0312, sig=0.531250)
x"3844", --  17  (x=0.0332, sig=0.533203)
x"3848", --  18  (x=0.0352, sig=0.535156)
x"384c", --  19  (x=0.0371, sig=0.537109)
x"3850", --  20  (x=0.0391, sig=0.539062)
x"3854", --  21  (x=0.0410, sig=0.541016)
x"3858", --  22  (x=0.0430, sig=0.542969)
x"385c", --  23  (x=0.0449, sig=0.544922)
x"3860", --  24  (x=0.0469, sig=0.546875)
x"3864", --  25  (x=0.0488, sig=0.548828)
x"3868", --  26  (x=0.0508, sig=0.550781)
x"386b", --  27  (x=0.0527, sig=0.552246)
x"386f", --  28  (x=0.0547, sig=0.554199)
x"3874", --  29  (x=0.0566, sig=0.556641)
x"3877", --  30  (x=0.0586, sig=0.558105)
x"387b", --  31  (x=0.0605, sig=0.560059)
x"387f", --  32  (x=0.0625, sig=0.562012)
x"3883", --  33  (x=0.0645, sig=0.563965)
x"3887", --  34  (x=0.0664, sig=0.565918)
x"388b", --  35  (x=0.0684, sig=0.567871)
x"388f", --  36  (x=0.0703, sig=0.569824)
x"3893", --  37  (x=0.0723, sig=0.571777)
x"3897", --  38  (x=0.0742, sig=0.573730)
x"389b", --  39  (x=0.0762, sig=0.575684)
x"389f", --  40  (x=0.0781, sig=0.577637)
x"38a2", --  41  (x=0.0801, sig=0.579102)
x"38a6", --  42  (x=0.0820, sig=0.581055)
x"38aa", --  43  (x=0.0840, sig=0.583008)
x"38ae", --  44  (x=0.0859, sig=0.584961)
x"38b2", --  45  (x=0.0879, sig=0.586914)
x"38b6", --  46  (x=0.0898, sig=0.588867)
x"38b9", --  47  (x=0.0918, sig=0.590332)
x"38be", --  48  (x=0.0938, sig=0.592773)
x"38c2", --  49  (x=0.0957, sig=0.594727)
x"38c5", --  50  (x=0.0977, sig=0.596191)
x"38c9", --  51  (x=0.0996, sig=0.598145)
x"38cd", --  52  (x=0.1016, sig=0.600098)
x"38d1", --  53  (x=0.1035, sig=0.602051)
x"38d5", --  54  (x=0.1055, sig=0.604004)
x"38d9", --  55  (x=0.1074, sig=0.605957)
x"38dd", --  56  (x=0.1094, sig=0.607910)
x"38e0", --  57  (x=0.1113, sig=0.609375)
x"38e4", --  58  (x=0.1133, sig=0.611328)
x"38e8", --  59  (x=0.1152, sig=0.613281)
x"38ec", --  60  (x=0.1172, sig=0.615234)
x"38ef", --  61  (x=0.1191, sig=0.616699)
x"38f3", --  62  (x=0.1211, sig=0.618652)
x"38f7", --  63  (x=0.1230, sig=0.620605)
x"38fb", --  64  (x=0.1250, sig=0.622559)
x"38ff", --  65  (x=0.1270, sig=0.624512)
x"3902", --  66  (x=0.1289, sig=0.625977)
x"3907", --  67  (x=0.1309, sig=0.628418)
x"390a", --  68  (x=0.1328, sig=0.629883)
x"390d", --  69  (x=0.1348, sig=0.631348)
x"3912", --  70  (x=0.1367, sig=0.633789)
x"3915", --  71  (x=0.1387, sig=0.635254)
x"3918", --  72  (x=0.1406, sig=0.636719)
x"391c", --  73  (x=0.1426, sig=0.638672)
x"3920", --  74  (x=0.1445, sig=0.640625)
x"3924", --  75  (x=0.1465, sig=0.642578)
x"3927", --  76  (x=0.1484, sig=0.644043)
x"392b", --  77  (x=0.1504, sig=0.645996)
x"392f", --  78  (x=0.1523, sig=0.647949)
x"3933", --  79  (x=0.1543, sig=0.649902)
x"3936", --  80  (x=0.1562, sig=0.651367)
x"3939", --  81  (x=0.1582, sig=0.652832)
x"393d", --  82  (x=0.1602, sig=0.654785)
x"3940", --  83  (x=0.1621, sig=0.656250)
x"3945", --  84  (x=0.1641, sig=0.658691)
x"3948", --  85  (x=0.1660, sig=0.660156)
x"394c", --  86  (x=0.1680, sig=0.662109)
x"394f", --  87  (x=0.1699, sig=0.663574)
x"3953", --  88  (x=0.1719, sig=0.665527)
x"3956", --  89  (x=0.1738, sig=0.666992)
x"395a", --  90  (x=0.1758, sig=0.668945)
x"395d", --  91  (x=0.1777, sig=0.670410)
x"3961", --  92  (x=0.1797, sig=0.672363)
x"3965", --  93  (x=0.1816, sig=0.674316)
x"3968", --  94  (x=0.1836, sig=0.675781)
x"396b", --  95  (x=0.1855, sig=0.677246)
x"396f", --  96  (x=0.1875, sig=0.679199)
x"3972", --  97  (x=0.1895, sig=0.680664)
x"3976", --  98  (x=0.1914, sig=0.682617)
x"397a", --  99  (x=0.1934, sig=0.684570)
x"397d", -- 100  (x=0.1953, sig=0.686035)
x"3980", -- 101  (x=0.1973, sig=0.687500)
x"3983", -- 102  (x=0.1992, sig=0.688965)
x"3987", -- 103  (x=0.2012, sig=0.690918)
x"398b", -- 104  (x=0.2031, sig=0.692871)
x"398e", -- 105  (x=0.2051, sig=0.694336)
x"3992", -- 106  (x=0.2070, sig=0.696289)
x"3995", -- 107  (x=0.2090, sig=0.697754)
x"3998", -- 108  (x=0.2109, sig=0.699219)
x"399b", -- 109  (x=0.2129, sig=0.700684)
x"399e", -- 110  (x=0.2148, sig=0.702148)
x"39a2", -- 111  (x=0.2168, sig=0.704102)
x"39a5", -- 112  (x=0.2188, sig=0.705566)
x"39a8", -- 113  (x=0.2207, sig=0.707031)
x"39ac", -- 114  (x=0.2227, sig=0.708984)
x"39af", -- 115  (x=0.2246, sig=0.710449)
x"39b2", -- 116  (x=0.2266, sig=0.711914)
x"39b6", -- 117  (x=0.2285, sig=0.713867)
x"39ba", -- 118  (x=0.2305, sig=0.715820)
x"39bd", -- 119  (x=0.2324, sig=0.717285)
x"39c0", -- 120  (x=0.2344, sig=0.718750)
x"39c3", -- 121  (x=0.2363, sig=0.720215)
x"39c6", -- 122  (x=0.2383, sig=0.721680)
x"39c9", -- 123  (x=0.2402, sig=0.723145)
x"39cc", -- 124  (x=0.2422, sig=0.724609)
x"39cf", -- 125  (x=0.2441, sig=0.726074)
x"39d3", -- 126  (x=0.2461, sig=0.728027)
x"39d6", -- 127  (x=0.2480, sig=0.729492)
x"39d9", -- 128  (x=0.2500, sig=0.730957)
x"39dc", -- 129  (x=0.2520, sig=0.732422)
x"39df", -- 130  (x=0.2539, sig=0.733887)
x"39e3", -- 131  (x=0.2559, sig=0.735840)
x"39e6", -- 132  (x=0.2578, sig=0.737305)
x"39e9", -- 133  (x=0.2598, sig=0.738770)
x"39eb", -- 134  (x=0.2617, sig=0.739746)
x"39ef", -- 135  (x=0.2637, sig=0.741699)
x"39f2", -- 136  (x=0.2656, sig=0.743164)
x"39f5", -- 137  (x=0.2676, sig=0.744629)
x"39f9", -- 138  (x=0.2695, sig=0.746582)
x"39fb", -- 139  (x=0.2715, sig=0.747559)
x"39fe", -- 140  (x=0.2734, sig=0.749023)
x"3a02", -- 141  (x=0.2754, sig=0.750977)
x"3a04", -- 142  (x=0.2773, sig=0.751953)
x"3a07", -- 143  (x=0.2793, sig=0.753418)
x"3a0b", -- 144  (x=0.2812, sig=0.755371)
x"3a0d", -- 145  (x=0.2832, sig=0.756348)
x"3a10", -- 146  (x=0.2852, sig=0.757812)
x"3a13", -- 147  (x=0.2871, sig=0.759277)
x"3a16", -- 148  (x=0.2891, sig=0.760742)
x"3a18", -- 149  (x=0.2910, sig=0.761719)
x"3a1c", -- 150  (x=0.2930, sig=0.763672)
x"3a1e", -- 151  (x=0.2949, sig=0.764648)
x"3a22", -- 152  (x=0.2969, sig=0.766602)
x"3a24", -- 153  (x=0.2988, sig=0.767578)
x"3a26", -- 154  (x=0.3008, sig=0.768555)
x"3a2a", -- 155  (x=0.3027, sig=0.770508)
x"3a2c", -- 156  (x=0.3047, sig=0.771484)
x"3a30", -- 157  (x=0.3066, sig=0.773438)
x"3a32", -- 158  (x=0.3086, sig=0.774414)
x"3a35", -- 159  (x=0.3105, sig=0.775879)
x"3a37", -- 160  (x=0.3125, sig=0.776855)
x"3a3b", -- 161  (x=0.3145, sig=0.778809)
x"3a3d", -- 162  (x=0.3164, sig=0.779785)
x"3a41", -- 163  (x=0.3184, sig=0.781738)
x"3a43", -- 164  (x=0.3203, sig=0.782715)
x"3a46", -- 165  (x=0.3223, sig=0.784180)
x"3a48", -- 166  (x=0.3242, sig=0.785156)
x"3a4b", -- 167  (x=0.3262, sig=0.786621)
x"3a4d", -- 168  (x=0.3281, sig=0.787598)
x"3a50", -- 169  (x=0.3301, sig=0.789062)
x"3a53", -- 170  (x=0.3320, sig=0.790527)
x"3a56", -- 171  (x=0.3340, sig=0.791992)
x"3a58", -- 172  (x=0.3359, sig=0.792969)
x"3a5b", -- 173  (x=0.3379, sig=0.794434)
x"3a5d", -- 174  (x=0.3398, sig=0.795410)
x"3a60", -- 175  (x=0.3418, sig=0.796875)
x"3a63", -- 176  (x=0.3438, sig=0.798340)
x"3a65", -- 177  (x=0.3457, sig=0.799316)
x"3a68", -- 178  (x=0.3477, sig=0.800781)
x"3a6a", -- 179  (x=0.3496, sig=0.801758)
x"3a6d", -- 180  (x=0.3516, sig=0.803223)
x"3a6f", -- 181  (x=0.3535, sig=0.804199)
x"3a72", -- 182  (x=0.3555, sig=0.805664)
x"3a75", -- 183  (x=0.3574, sig=0.807129)
x"3a77", -- 184  (x=0.3594, sig=0.808105)
x"3a7a", -- 185  (x=0.3613, sig=0.809570)
x"3a7b", -- 186  (x=0.3633, sig=0.810059)
x"3a7e", -- 187  (x=0.3652, sig=0.811523)
x"3a80", -- 188  (x=0.3672, sig=0.812500)
x"3a83", -- 189  (x=0.3691, sig=0.813965)
x"3a86", -- 190  (x=0.3711, sig=0.815430)
x"3a88", -- 191  (x=0.3730, sig=0.816406)
x"3a8b", -- 192  (x=0.3750, sig=0.817871)
x"3a8c", -- 193  (x=0.3770, sig=0.818359)
x"3a8f", -- 194  (x=0.3789, sig=0.819824)
x"3a92", -- 195  (x=0.3809, sig=0.821289)
x"3a93", -- 196  (x=0.3828, sig=0.821777)
x"3a96", -- 197  (x=0.3848, sig=0.823242)
x"3a99", -- 198  (x=0.3867, sig=0.824707)
x"3a9b", -- 199  (x=0.3887, sig=0.825684)
x"3a9d", -- 200  (x=0.3906, sig=0.826660)
x"3a9f", -- 201  (x=0.3926, sig=0.827637)
x"3aa2", -- 202  (x=0.3945, sig=0.829102)
x"3aa3", -- 203  (x=0.3965, sig=0.829590)
x"3aa6", -- 204  (x=0.3984, sig=0.831055)
x"3aa9", -- 205  (x=0.4004, sig=0.832520)
x"3aaa", -- 206  (x=0.4023, sig=0.833008)
x"3aad", -- 207  (x=0.4043, sig=0.834473)
x"3aaf", -- 208  (x=0.4062, sig=0.835449)
x"3ab1", -- 209  (x=0.4082, sig=0.836426)
x"3ab4", -- 210  (x=0.4102, sig=0.837891)
x"3ab6", -- 211  (x=0.4121, sig=0.838867)
x"3ab8", -- 212  (x=0.4141, sig=0.839844)
x"3aba", -- 213  (x=0.4160, sig=0.840820)
x"3abd", -- 214  (x=0.4180, sig=0.842285)
x"3abe", -- 215  (x=0.4199, sig=0.842773)
x"3ac1", -- 216  (x=0.4219, sig=0.844238)
x"3ac2", -- 217  (x=0.4238, sig=0.844727)
x"3ac5", -- 218  (x=0.4258, sig=0.846191)
x"3ac7", -- 219  (x=0.4277, sig=0.847168)
x"3ac8", -- 220  (x=0.4297, sig=0.847656)
x"3acb", -- 221  (x=0.4316, sig=0.849121)
x"3acc", -- 222  (x=0.4336, sig=0.849609)
x"3acf", -- 223  (x=0.4355, sig=0.851074)
x"3ad1", -- 224  (x=0.4375, sig=0.852051)
x"3ad4", -- 225  (x=0.4395, sig=0.853516)
x"3ad5", -- 226  (x=0.4414, sig=0.854004)
x"3ad7", -- 227  (x=0.4434, sig=0.854980)
x"3ad9", -- 228  (x=0.4453, sig=0.855957)
x"3adb", -- 229  (x=0.4473, sig=0.856934)
x"3adc", -- 230  (x=0.4492, sig=0.857422)
x"3adf", -- 231  (x=0.4512, sig=0.858887)
x"3ae1", -- 232  (x=0.4531, sig=0.859863)
x"3ae2", -- 233  (x=0.4551, sig=0.860352)
x"3ae4", -- 234  (x=0.4570, sig=0.861328)
x"3ae7", -- 235  (x=0.4590, sig=0.862793)
x"3ae8", -- 236  (x=0.4609, sig=0.863281)
x"3aea", -- 237  (x=0.4629, sig=0.864258)
x"3aeb", -- 238  (x=0.4648, sig=0.864746)
x"3aee", -- 239  (x=0.4668, sig=0.866211)
x"3af0", -- 240  (x=0.4688, sig=0.867188)
x"3af1", -- 241  (x=0.4707, sig=0.867676)
x"3af3", -- 242  (x=0.4727, sig=0.868652)
x"3af6", -- 243  (x=0.4746, sig=0.870117)
x"3af7", -- 244  (x=0.4766, sig=0.870605)
x"3af9", -- 245  (x=0.4785, sig=0.871582)
x"3afa", -- 246  (x=0.4805, sig=0.872070)
x"3afc", -- 247  (x=0.4824, sig=0.873047)
x"3afd", -- 248  (x=0.4844, sig=0.873535)
x"3b00", -- 249  (x=0.4863, sig=0.875000)
x"3b02", -- 250  (x=0.4883, sig=0.875977)
x"3b04", -- 251  (x=0.4902, sig=0.876953)
x"3b05", -- 252  (x=0.4922, sig=0.877441)
x"3b07", -- 253  (x=0.4941, sig=0.878418)
x"3b08", -- 254  (x=0.4961, sig=0.878906)
x"3b0a", -- 255  (x=0.4980, sig=0.879883)
x"3b0b", -- 256  (x=0.5000, sig=0.880371)
x"3b10", -- 257  (x=0.5039, sig=0.882812)
x"3b13", -- 258  (x=0.5078, sig=0.884277)
x"3b16", -- 259  (x=0.5117, sig=0.885742)
x"3b19", -- 260  (x=0.5156, sig=0.887207)
x"3b1c", -- 261  (x=0.5195, sig=0.888672)
x"3b20", -- 262  (x=0.5234, sig=0.890625)
x"3b23", -- 263  (x=0.5273, sig=0.892090)
x"3b26", -- 264  (x=0.5312, sig=0.893555)
x"3b29", -- 265  (x=0.5352, sig=0.895020)
x"3b2b", -- 266  (x=0.5391, sig=0.895996)
x"3b2e", -- 267  (x=0.5430, sig=0.897461)
x"3b31", -- 268  (x=0.5469, sig=0.898926)
x"3b34", -- 269  (x=0.5508, sig=0.900391)
x"3b38", -- 270  (x=0.5547, sig=0.902344)
x"3b39", -- 271  (x=0.5586, sig=0.902832)
x"3b3d", -- 272  (x=0.5625, sig=0.904785)
x"3b40", -- 273  (x=0.5664, sig=0.906250)
x"3b42", -- 274  (x=0.5703, sig=0.907227)
x"3b45", -- 275  (x=0.5742, sig=0.908691)
x"3b48", -- 276  (x=0.5781, sig=0.910156)
x"3b4a", -- 277  (x=0.5820, sig=0.911133)
x"3b4d", -- 278  (x=0.5859, sig=0.912598)
x"3b4f", -- 279  (x=0.5898, sig=0.913574)
x"3b52", -- 280  (x=0.5938, sig=0.915039)
x"3b54", -- 281  (x=0.5977, sig=0.916016)
x"3b57", -- 282  (x=0.6016, sig=0.917480)
x"3b59", -- 283  (x=0.6055, sig=0.918457)
x"3b5b", -- 284  (x=0.6094, sig=0.919434)
x"3b5e", -- 285  (x=0.6133, sig=0.920898)
x"3b60", -- 286  (x=0.6172, sig=0.921875)
x"3b63", -- 287  (x=0.6211, sig=0.923340)
x"3b65", -- 288  (x=0.6250, sig=0.924316)
x"3b66", -- 289  (x=0.6289, sig=0.924805)
x"3b68", -- 290  (x=0.6328, sig=0.925781)
x"3b6c", -- 291  (x=0.6367, sig=0.927734)
x"3b6d", -- 292  (x=0.6406, sig=0.928223)
x"3b6f", -- 293  (x=0.6445, sig=0.929199)
x"3b71", -- 294  (x=0.6484, sig=0.930176)
x"3b74", -- 295  (x=0.6523, sig=0.931641)
x"3b76", -- 296  (x=0.6562, sig=0.932617)
x"3b78", -- 297  (x=0.6602, sig=0.933594)
x"3b79", -- 298  (x=0.6641, sig=0.934082)
x"3b7b", -- 299  (x=0.6680, sig=0.935059)
x"3b7d", -- 300  (x=0.6719, sig=0.936035)
x"3b7f", -- 301  (x=0.6758, sig=0.937012)
x"3b80", -- 302  (x=0.6797, sig=0.937500)
x"3b84", -- 303  (x=0.6836, sig=0.939453)
x"3b86", -- 304  (x=0.6875, sig=0.940430)
x"3b88", -- 305  (x=0.6914, sig=0.941406)
x"3b89", -- 306  (x=0.6953, sig=0.941895)
x"3b8b", -- 307  (x=0.6992, sig=0.942871)
x"3b8b", -- 308  (x=0.7031, sig=0.942871)
x"3b8d", -- 309  (x=0.7070, sig=0.943848)
x"3b8f", -- 310  (x=0.7109, sig=0.944824)
x"3b90", -- 311  (x=0.7148, sig=0.945312)
x"3b92", -- 312  (x=0.7188, sig=0.946289)
x"3b94", -- 313  (x=0.7227, sig=0.947266)
x"3b96", -- 314  (x=0.7266, sig=0.948242)
x"3b98", -- 315  (x=0.7305, sig=0.949219)
x"3b99", -- 316  (x=0.7344, sig=0.949707)
x"3b9b", -- 317  (x=0.7383, sig=0.950684)
x"3b9b", -- 318  (x=0.7422, sig=0.950684)
x"3b9d", -- 319  (x=0.7461, sig=0.951660)
x"3b9f", -- 320  (x=0.7500, sig=0.952637)
x"3ba1", -- 321  (x=0.7539, sig=0.953613)
x"3ba2", -- 322  (x=0.7578, sig=0.954102)
x"3ba2", -- 323  (x=0.7617, sig=0.954102)
x"3ba4", -- 324  (x=0.7656, sig=0.955078)
x"3ba6", -- 325  (x=0.7695, sig=0.956055)
x"3ba8", -- 326  (x=0.7734, sig=0.957031)
x"3ba8", -- 327  (x=0.7773, sig=0.957031)
x"3baa", -- 328  (x=0.7812, sig=0.958008)
x"3bac", -- 329  (x=0.7852, sig=0.958984)
x"3bac", -- 330  (x=0.7891, sig=0.958984)
x"3bad", -- 331  (x=0.7930, sig=0.959473)
x"3baf", -- 332  (x=0.7969, sig=0.960449)
x"3baf", -- 333  (x=0.8008, sig=0.960449)
x"3bb1", -- 334  (x=0.8047, sig=0.961426)
x"3bb3", -- 335  (x=0.8086, sig=0.962402)
x"3bb3", -- 336  (x=0.8125, sig=0.962402)
x"3bb5", -- 337  (x=0.8164, sig=0.963379)
x"3bb7", -- 338  (x=0.8203, sig=0.964355)
x"3bb7", -- 339  (x=0.8242, sig=0.964355)
x"3bb9", -- 340  (x=0.8281, sig=0.965332)
x"3bb9", -- 341  (x=0.8320, sig=0.965332)
x"3bba", -- 342  (x=0.8359, sig=0.965820)
x"3bba", -- 343  (x=0.8398, sig=0.965820)
x"3bbc", -- 344  (x=0.8438, sig=0.966797)
x"3bbe", -- 345  (x=0.8477, sig=0.967773)
x"3bbe", -- 346  (x=0.8516, sig=0.967773)
x"3bc0", -- 347  (x=0.8555, sig=0.968750)
x"3bc0", -- 348  (x=0.8594, sig=0.968750)
x"3bc2", -- 349  (x=0.8633, sig=0.969727)
x"3bc2", -- 350  (x=0.8672, sig=0.969727)
x"3bc4", -- 351  (x=0.8711, sig=0.970703)
x"3bc4", -- 352  (x=0.8750, sig=0.970703)
x"3bc6", -- 353  (x=0.8789, sig=0.971680)
x"3bc6", -- 354  (x=0.8828, sig=0.971680)
x"3bc6", -- 355  (x=0.8867, sig=0.971680)
x"3bc8", -- 356  (x=0.8906, sig=0.972656)
x"3bc8", -- 357  (x=0.8945, sig=0.972656)
x"3bc9", -- 358  (x=0.8984, sig=0.973145)
x"3bc9", -- 359  (x=0.9023, sig=0.973145)
x"3bcb", -- 360  (x=0.9062, sig=0.974121)
x"3bcb", -- 361  (x=0.9102, sig=0.974121)
x"3bcd", -- 362  (x=0.9141, sig=0.975098)
x"3bcd", -- 363  (x=0.9180, sig=0.975098)
x"3bcd", -- 364  (x=0.9219, sig=0.975098)
x"3bcf", -- 365  (x=0.9258, sig=0.976074)
x"3bcf", -- 366  (x=0.9297, sig=0.976074)
x"3bd1", -- 367  (x=0.9336, sig=0.977051)
x"3bd1", -- 368  (x=0.9375, sig=0.977051)
x"3bd1", -- 369  (x=0.9414, sig=0.977051)
x"3bd3", -- 370  (x=0.9453, sig=0.978027)
x"3bd3", -- 371  (x=0.9492, sig=0.978027)
x"3bd3", -- 372  (x=0.9531, sig=0.978027)
x"3bd5", -- 373  (x=0.9570, sig=0.979004)
x"3bd5", -- 374  (x=0.9609, sig=0.979004)
x"3bd5", -- 375  (x=0.9648, sig=0.979004)
x"3bd7", -- 376  (x=0.9688, sig=0.979980)
x"3bd7", -- 377  (x=0.9727, sig=0.979980)
x"3bd7", -- 378  (x=0.9766, sig=0.979980)
x"3bd9", -- 379  (x=0.9805, sig=0.980957)
x"3bd9", -- 380  (x=0.9844, sig=0.980957)
x"3bd9", -- 381  (x=0.9883, sig=0.980957)
x"3bdb", -- 382  (x=0.9922, sig=0.981934)
x"3bdb", -- 383  (x=0.9961, sig=0.981934)
x"3bdb", -- 384  (x=1.0000, sig=0.981934)
x"3bdd", -- 385  (x=1.0078, sig=0.982910)
x"3bdd", -- 386  (x=1.0156, sig=0.982910)
x"3bdf", -- 387  (x=1.0234, sig=0.983887)
x"3bdf", -- 388  (x=1.0312, sig=0.983887)
x"3be0", -- 389  (x=1.0391, sig=0.984375)
x"3be0", -- 390  (x=1.0469, sig=0.984375)
x"3be2", -- 391  (x=1.0547, sig=0.985352)
x"3be2", -- 392  (x=1.0625, sig=0.985352)
x"3be4", -- 393  (x=1.0703, sig=0.986328)
x"3be4", -- 394  (x=1.0781, sig=0.986328)
x"3be6", -- 395  (x=1.0859, sig=0.987305)
x"3be6", -- 396  (x=1.0938, sig=0.987305)
x"3be8", -- 397  (x=1.1016, sig=0.988281)
x"3be8", -- 398  (x=1.1094, sig=0.988281)
x"3be8", -- 399  (x=1.1172, sig=0.988281)
x"3bea", -- 400  (x=1.1250, sig=0.989258)
x"3bea", -- 401  (x=1.1328, sig=0.989258)
x"3bea", -- 402  (x=1.1406, sig=0.989258)
x"3bec", -- 403  (x=1.1484, sig=0.990234)
x"3bec", -- 404  (x=1.1562, sig=0.990234)
x"3bec", -- 405  (x=1.1641, sig=0.990234)
x"3bee", -- 406  (x=1.1719, sig=0.991211)
x"3bee", -- 407  (x=1.1797, sig=0.991211)
x"3bee", -- 408  (x=1.1875, sig=0.991211)
x"3bee", -- 409  (x=1.1953, sig=0.991211)
x"3bf0", -- 410  (x=1.2031, sig=0.992188)
x"3bf0", -- 411  (x=1.2109, sig=0.992188)
x"3bf0", -- 412  (x=1.2188, sig=0.992188)
x"3bf0", -- 413  (x=1.2266, sig=0.992188)
x"3bf2", -- 414  (x=1.2344, sig=0.993164)
x"3bf2", -- 415  (x=1.2422, sig=0.993164)
x"3bf2", -- 416  (x=1.2500, sig=0.993164)
x"3bf2", -- 417  (x=1.2578, sig=0.993164)
x"3bf4", -- 418  (x=1.2656, sig=0.994141)
x"3bf4", -- 419  (x=1.2734, sig=0.994141)
x"3bf4", -- 420  (x=1.2812, sig=0.994141)
x"3bf4", -- 421  (x=1.2891, sig=0.994141)
x"3bf4", -- 422  (x=1.2969, sig=0.994141)
x"3bf4", -- 423  (x=1.3047, sig=0.994141)
x"3bf6", -- 424  (x=1.3125, sig=0.995117)
x"3bf6", -- 425  (x=1.3203, sig=0.995117)
x"3bf6", -- 426  (x=1.3281, sig=0.995117)
x"3bf6", -- 427  (x=1.3359, sig=0.995117)
x"3bf6", -- 428  (x=1.3438, sig=0.995117)
x"3bf6", -- 429  (x=1.3516, sig=0.995117)
x"3bf8", -- 430  (x=1.3594, sig=0.996094)
x"3bf8", -- 431  (x=1.3672, sig=0.996094)
x"3bf8", -- 432  (x=1.3750, sig=0.996094)
x"3bf8", -- 433  (x=1.3828, sig=0.996094)
x"3bf8", -- 434  (x=1.3906, sig=0.996094)
x"3bf8", -- 435  (x=1.3984, sig=0.996094)
x"3bf8", -- 436  (x=1.4062, sig=0.996094)
x"3bf8", -- 437  (x=1.4141, sig=0.996094)
x"3bfa", -- 438  (x=1.4219, sig=0.997070)
x"3bfa", -- 439  (x=1.4297, sig=0.997070)
x"3bfa", -- 440  (x=1.4375, sig=0.997070)
x"3bfa", -- 441  (x=1.4453, sig=0.997070)
x"3bfa", -- 442  (x=1.4531, sig=0.997070)
x"3bfa", -- 443  (x=1.4609, sig=0.997070)
x"3bfa", -- 444  (x=1.4688, sig=0.997070)
x"3bfa", -- 445  (x=1.4766, sig=0.997070)
x"3bfa", -- 446  (x=1.4844, sig=0.997070)
x"3bfa", -- 447  (x=1.4922, sig=0.997070)
x"3bfa", -- 448  (x=1.5000, sig=0.997070)
x"3bfc", -- 449  (x=1.5078, sig=0.998047)
x"3bfc", -- 450  (x=1.5156, sig=0.998047)
x"3bfc", -- 451  (x=1.5234, sig=0.998047)
x"3bfc", -- 452  (x=1.5312, sig=0.998047)
x"3bfc", -- 453  (x=1.5400, sig=0.998047)
x"3bfc", -- 454  (x=1.5479, sig=0.998047)
x"3bfc", -- 455  (x=1.5557, sig=0.998047)
x"3bfc", -- 456  (x=1.5635, sig=0.998047)
x"3bfc", -- 457  (x=1.5713, sig=0.998047)
x"3bfc", -- 458  (x=1.5791, sig=0.998047)
x"3bfc", -- 459  (x=1.5869, sig=0.998047)
x"3bfc", -- 460  (x=1.5957, sig=0.998047)
x"3bfc", -- 461  (x=1.6035, sig=0.998047)
x"3bfc", -- 462  (x=1.6113, sig=0.998047)
x"3bfc", -- 463  (x=1.6191, sig=0.998047)
x"3bfc", -- 464  (x=1.6270, sig=0.998047)
x"3bfe", -- 465  (x=1.6348, sig=0.999023)
x"3bfe", -- 466  (x=1.6426, sig=0.999023)
x"3bfe", -- 467  (x=1.6504, sig=0.999023)
x"3bfe", -- 468  (x=1.6582, sig=0.999023)
x"3bfe", -- 469  (x=1.6670, sig=0.999023)
x"3bfe", -- 470  (x=1.6748, sig=0.999023)
x"3bfe", -- 471  (x=1.6826, sig=0.999023)
x"3bfe", -- 472  (x=1.6904, sig=0.999023)
x"3bfe", -- 473  (x=1.6982, sig=0.999023)
x"3bfe", -- 474  (x=1.7061, sig=0.999023)
x"3bfe", -- 475  (x=1.7139, sig=0.999023)
x"3bfe", -- 476  (x=1.7227, sig=0.999023)
x"3bfe", -- 477  (x=1.7305, sig=0.999023)
x"3bfe", -- 478  (x=1.7383, sig=0.999023)
x"3bfe", -- 479  (x=1.7461, sig=0.999023)
x"3bfe", -- 480  (x=1.7539, sig=0.999023)
x"3bfe", -- 481  (x=1.7617, sig=0.999023)
x"3bfe", -- 482  (x=1.7695, sig=0.999023)
x"3bfe", -- 483  (x=1.7773, sig=0.999023)
x"3bfe", -- 484  (x=1.7852, sig=0.999023)
x"3bfe", -- 485  (x=1.7930, sig=0.999023)
x"3bfe", -- 486  (x=1.8018, sig=0.999023)
x"3bfe", -- 487  (x=1.8096, sig=0.999023)
x"3bfe", -- 488  (x=1.8174, sig=0.999023)
x"3bfe", -- 489  (x=1.8252, sig=0.999023)
x"3bfe", -- 490  (x=1.8330, sig=0.999023)
x"3bfe", -- 491  (x=1.8418, sig=0.999023)
x"3bfe", -- 492  (x=1.8496, sig=0.999023)
x"3bfe", -- 493  (x=1.8574, sig=0.999023)
x"3bfe", -- 494  (x=1.8652, sig=0.999023)
x"3bfe", -- 495  (x=1.8730, sig=0.999023)
x"3bfe", -- 496  (x=1.8809, sig=0.999023)
x"3bfe", -- 497  (x=1.8887, sig=0.999023)
x"3bfe", -- 498  (x=1.8965, sig=0.999023)
x"3bfe", -- 499  (x=1.9043, sig=0.999023)
x"3c00", -- 500  (x=1.9121, sig=1.000000)
x"3c00", -- 501  (x=1.9199, sig=1.000000)
x"3c00", -- 502  (x=1.9287, sig=1.000000)
x"3c00", -- 503  (x=1.9365, sig=1.000000)
x"3c00", -- 504  (x=1.9443, sig=1.000000)
x"3c00", -- 505  (x=1.9521, sig=1.000000)
x"3c00", -- 506  (x=1.9600, sig=1.000000)
x"3c00", -- 507  (x=1.9688, sig=1.000000)
x"3c00", -- 508  (x=1.9766, sig=1.000000)
x"3c00", -- 509  (x=1.9844, sig=1.000000)
x"3c00", -- 510  (x=1.9922, sig=1.000000)
x"3c00" -- 511  (x=2.0000, sig=1.000000)


    );
end package LUT;


